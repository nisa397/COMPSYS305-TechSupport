library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_lfsr is
end entity tb_lfsr;

architecture arc of tb_lfsr is

	component lfsr
		port( seed: in unsigned(7 downto 0);
		Clock: in std_logic;
		rand_num: out unsigned(7 downto 0));  
	end component;
	
	signal Clk_tb: std_logic := '0';
	signal seed_tb: unsigned (7 downto 0) := to_unsigned(114, 8);
	signal rand_tb: unsigned (7 downto 0);
begin
	
	LFSR_TB:lfsr 
	port map(
	seed => seed_tb,
	Clock => Clk_tb,
	rand_num => rand_tb
	);

	process
	begin
	CLK_tb <= '0';
   	wait for 5 ns;
    	CLK_tb <= '1';
    	wait for 5 ns;
	end process;
end arc;

	
	
